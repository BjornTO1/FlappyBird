module rand_pipe (random, pipe);
input logic [3:0] random;
output logic [15:0][15:0] pipe;

always_comb begin 
	casex(random)
		4'b1xxx: begin pipe[00] = 16'b0000000000000001;
					pipe[01] = 16'b0000000000000000;
					pipe[02] = 16'b0000000000000000;
					pipe[03] = 16'b0000000000000000;
					pipe[04] = 16'b0000000000000000;
					pipe[05] = 16'b0000000000000001;
					pipe[06] = 16'b0000000000000001;
					pipe[07] = 16'b0000000000000001;
					pipe[08] = 16'b0000000000000001;
					pipe[09] = 16'b0000000000000001;
					pipe[10] = 16'b0000000000000001;
					pipe[11] = 16'b0000000000000001;
					pipe[12] = 16'b0000000000000001;
					pipe[13] = 16'b0000000000000001;
					pipe[14] = 16'b0000000000000001;
					pipe[15] = 16'b0000000000000001;
					end
							 
		4'b01xx: begin pipe[00] = 16'b0000000000000001;
					pipe[01] = 16'b0000000000000001;
					pipe[02] = 16'b0000000000000001;
					pipe[03] = 16'b0000000000000001;
					pipe[04] = 16'b0000000000000000;
					pipe[05] = 16'b0000000000000000;
					pipe[06] = 16'b0000000000000000;
				   pipe[07] = 16'b0000000000000000;
					pipe[08] = 16'b0000000000000001;
					pipe[09] = 16'b0000000000000001;
					pipe[10] = 16'b0000000000000001;
					pipe[11] = 16'b0000000000000001;
					pipe[12] = 16'b0000000000000001;
					pipe[13] = 16'b0000000000000001;
					pipe[14] = 16'b0000000000000001;
					pipe[15] = 16'b0000000000000001;
					end
					
		4'b001x: begin pipe[00] = 16'b0000000000000001;
					pipe[01] = 16'b0000000000000001;
					pipe[02] = 16'b0000000000000001;
					pipe[03] = 16'b0000000000000001;
					pipe[04] = 16'b0000000000000001;
					pipe[05] = 16'b0000000000000001;
					pipe[06] = 16'b0000000000000001;
				   pipe[07] = 16'b0000000000000001;
					pipe[08] = 16'b0000000000000000;
					pipe[09] = 16'b0000000000000000;
					pipe[10] = 16'b0000000000000000;
					pipe[11] = 16'b0000000000000000;
					pipe[12] = 16'b0000000000000001;
					pipe[13] = 16'b0000000000000001;
					pipe[14] = 16'b0000000000000001;
					pipe[15] = 16'b0000000000000001;
					end
					
		4'b0001: begin pipe[00] = 16'b0000000000000001;
					pipe[01] = 16'b0000000000000001;
					pipe[02] = 16'b0000000000000001;
					pipe[03] = 16'b0000000000000001;
					pipe[04] = 16'b0000000000000001;
					pipe[05] = 16'b0000000000000001;
					pipe[06] = 16'b0000000000000001;
				   pipe[07] = 16'b0000000000000001;
					pipe[08] = 16'b0000000000000001;
					pipe[09] = 16'b0000000000000001;
					pipe[10] = 16'b0000000000000001;
					pipe[11] = 16'b0000000000000000;
					pipe[12] = 16'b0000000000000000;
					pipe[13] = 16'b0000000000000000;
					pipe[14] = 16'b0000000000000000;
					pipe[15] = 16'b0000000000000001;
					end
	endcase
end

endmodule
